`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2024/05/08 20:37:20
// Design Name: 
// Module Name: insmem
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module insmem(addr_code, code);
input [5:0] addr_code;
output reg [31:0] code;

reg [31:0] mem [63:0];
initial begin
//flow water test code�� which is used for verifying I-type code
      mem[0] = 32'b10000000_00000000_00000100_000010_01;
      mem[1] = 32'b10000000_00000001_00000101_000011_01;
      mem[2] = 32'b01000000_00000001_00000110_000011_01;
      mem[3] = 32'b00100000_00000001_00000111_000011_01;
      mem[4] = 32'b00010000_00000001_00001000_000011_01;
      mem[5] = 32'b00001000_00000001_00001001_000011_01;
      mem[6] = 32'b00000100_00000001_00001010_000011_01;
      mem[7] = 32'b00000010_00000001_00001011_000011_01;

//load, store, move test code
//        mem[0] = 32'b00000000_00000001_00001000_000000_10;      
//          mem[0] = 32'b00000000_00001000_00000000_000001_10;
//          mem[1] = 32'b00000000_00000001_00001000_000000_10;
//          mem[2] = 32'b00000000_00000001_00001000_000010_10;

//verification of R,I tupe code
//        mem[0] = 32'b00000000_00000001_00001001_000000_00;
//        mem[1] = 32'b00000000_00000001_00001001_000001_00;
//        mem[2] = 32'b00000011_00000000_00001001_000000_01;
//        mem[3] = 32'b00000011_00000000_00001011_000001_01;



//        mem[1] = 32'b00000000_10000001_00000001_000001_10;
//        mem[2] = 32'b00000000_00000001_10000000_000010_10;
//      mem[8] = 32'b00000000_00000111_00000001_000000_10;
//      mem[9] = 32'b00000000_00000001_00000111_000001_10;
//      mem[10] = 32'b00000000_00000001_00000011_000010_10;
//    mem[0] = 32'b00000010_00000000_00000010_000010_01;
//    mem[1] = 32'b00000010_00000010_00000011_000010_01;
//    mem[2] = 32'b00000010_00000011_00000100_000010_01;
//    mem[3] = 32'b00000010_00000100_00000101_000010_01;
//    mem[4] = 32'b00000010_00000101_00000110_000010_01;
//    mem[5] = 32'b00000010_00000110_00000111_000010_01;
//    mem[6] = 32'b00000010_00000111_00001000_000010_01;
//    mem[7] = 32'b00000010_00000111_00001000_000010_01;
//mem[4] = 32'b00000000_00000001_00000010_000010_00;
//mem[6] = 32'b00000000_00000001_00000010_000011_00;
//mem[8] = 32'b00000000_00000001_00000010_000100_00;
//mem[10] = 32'b00000000_00000001_00000010_000101_00;
//mem[12] = 32'b00000000_00000001_00000010_000110_00;
//mem[14] = 32'b00000000_00000001_00000010_000111_00;
//mem[16] = 32'b00000000_00000001_00000010_001000_00;
//mem[18] = 32'b00000000_00000001_00000010_001001_00;
//mem[20] = 32'b00000000_00000001_00000010_001010_00;
//mem[22] = 32'b00000000_00000001_00000010_001011_00;
//mem[24] = 32'b00000000_00000001_00000010_001100_00;
//  mem[2] = 32'b00000011_00000001_00000010_000000_01;//26
//  mem[3] = 32'b00000011_00000001_00000010_000001_01;//30
//mem[32] = 32'b00000011_00000001_00000010_000010_01;
//mem[34] = 32'b00000011_00000001_00000010_000011_01;
//mem[36] = 32'b00000011_00000001_00000010_000100_01;
//mem[38] = 32'b00000011_00000001_00000010_000101_01;
//mem[40] = 32'b00000011_00000001_00000010_000110_01;
//mem[42] = 32'b00000011_00000001_00000010_000111_01;
//mem[44] = 32'b00000011_00000001_00000010_001000_01;
//mem[46] = 32'b00000011_00000001_00000010_001001_01;
//mem[48] = 32'b00000011_00000001_00000010_001010_01;
//mem[50] = 32'b00000011_00000001_00000010_001011_01;
//mem[52] = 32'b00000011_00000001_00000010_001100_01;
//mem[4] = 32'b00000000_00000001_00010000_000000_10;//54
//mem[5] = 32'b00000000_00010000_00000000_000001_10;//56
//mem[6] = 32'b00000000_00000001_00010000_000010_10;//58
end
always@(*)
begin
  code = mem[addr_code];
end
endmodule
